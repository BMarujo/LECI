library IEEE;
use IEEE.STD_LOGIC_1164.all;

-- Entidade sem portos
entity CounterUpDown_Tb is
end CounterUpDown_Tb;

architecture Stimulus of CounterUpDown_Tb is
 -- Sinais para ligar às entradas da UUT
	signal s_reset, s_clk : std_logic;
	signal s_upDown_n : std_logic;

 -- Sinal para ligar às saídas da UUT
	signal s_cntOut : std_logic_vector(3 downto 0);
begin
 -- Instanciação da Unit Under Test (UUT)
	uut : entity work.CounterUpDown4(Behavioral)
			port map(reset => s_reset,
						clk => s_clk,
						upDown => s_upDown_n,
						count => s_cntOut);
						
 -- Process clock
	 clock_proc : process
	 begin
		s_clk <= '0'; wait for 100 ns;
		s_clk <= '1'; wait for 100 ns;
	end process;

 --Process stim
 stim_proc : process
 begin
		s_reset <= '1';
		s_upDown_n <= '1';
		wait for 325 ns;
		s_reset <= '0';
		wait for 325 ns;
		s_upDown_n <= '0';
		wait for 325 ns;
		s_reset <= '1';
		wait for 325 ns;
		s_reset <= '0';
		s_upDown_n <= '1';
		wait for 950 ns;
	end process;
end Stimulus; 