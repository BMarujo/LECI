library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Machine is
	port(reset : in std_logic;
		  clk : in std_logic;
		  input : in std_logic_vector(1 downto 0);
		  output : out std_logic);
end Machine;

architecture Behavioral of Machine is
	type TState is (S0,S1,S2,S3,S4,S5);
	signal pState, nState: TState;
	
begin
	sync_proc : process(clk)
	begin
		if (rising_edge(clk)) then
			if (reset = '1') then
				pState <= S0;
			else
				pState <= nState;
			end if;
		end if;
end process;

	comb_proc : process(pState, input)
	begin
		case pState is
			when S0 =>
				output <= '0'; -- Moore output
				if (input(0) = '1') then
					nState <= S1;
				elsif(input(1) = '1') then
					nState <= S3;
				end if;
					
			when S1 =>
				output <= '0'; -- Moore output
				if (input(0) = '1') then
					nState <= S2;
				elsif(input(1) = '1') then
					nState <= S4;
				end if;
					
			when S2 =>
				output <= '0'; -- Moore output
				if (input(0) = '1') then
					nState <= S3;
				elsif(input(1) = '1') then
					nState <= S5;
				end if;
					
			when S3 =>
				output <= '0'; -- Moore output
				if (input(0) = '1') then
					nState <= S4;
				elsif(input(1) = '1') then
					nState <= S5;
				end if;
					
			when S4 =>
				output <= '0'; -- Moore output
				if (input(0) = '1' or input(1) = '1') then
					nState <= S5;
				end if;
				
			when S5 =>
				output <= '1';
				nState <= S0;
				
			when others => -- “Catch all” condition
					nState <= S0;
					output <= '0';
		end case;
	end process;
end Behavioral;