library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity CombShiftUnit_Demo is
	port(CLOCK_50 : in std_logic;
		  SW  : in std_logic_vector(10 downto 0);
		  KEY : in std_logic_vector(2 downto 0);
		  LEDR: out std_logic_vector(7 downto 0));
end CombShiftUnit_Demo;
architecture Behavioral of CombShiftUnit_Demo is
	signal clkout : std_logic;
begin
	clocky: entity work.ClkDividerN(Behavioral)
			  generic map(divFactor => 50000000) 
			  port map(clkIn => CLOCK_50,
						  clkOut => clkout);
	
	Combo : entity work.CombShiftUnit(Behavioral)
			  port map(clk=>clkout,
						  dataIn=>SW(7 downto 0),
						  rotate=>KEY(0),
						  dirLeft=>KEY(1),
						  shArith=>KEY(2),
						  shAmount=>SW(10 downto 8),
						  dataOut=>LEDR(7 downto 0));
end Behavioral;